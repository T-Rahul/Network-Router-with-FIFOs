  module router_fsm (clock, resetn, pkt_valid, data_in, fifo_full, fifo_empty_0, fifo_empty_1, fifo_empty_2, soft_reset_0, soft_reset_1, soft_reset_2, parity_done, low_packet_valid,
                     write_enb_reg, detect_add, ld_state, laf_state, lfd_state, full_state, rst_int_reg, busy);
  
  input clock, resetn, pkt_valid, fifo_full, fifo_empty_0, fifo_empty_1, fifo_empty_2, soft_reset_0, soft_reset_1, soft_reset_2, parity_done, low_packet_valid;
  input [1:0] data_in;
  output write_enb_reg, detect_add, ld_state, laf_state, lfd_state, full_state, rst_int_reg, busy;
  
  parameter DA  = 3'd0;  //DECODE_ADDRESS
  parameter LFD = 3'd1;  //LOAD_FIRST_DATA
  parameter LD  = 3'd2;  //LOAD_DATA
  parameter LP  = 3'd3;  //LOAD_PARITY
  parameter FFS = 3'd4;  //FIFO_FULL_STATE
  parameter LAF = 3'd5;  //LOAD_AFTER_FULL
  parameter WTE = 3'd6;  //WAIT_TILL_EMPTY
  parameter CPE = 3'd7;  //CHECK_PARITY_ERROR
  
  reg [2:0] state, next_state;
  
  always@(posedge clock, negedge resetn)
  begin
  
  if(!resetn)
  state <= DA;
  else if(((data_in == 2'b00) && soft_reset_0) ||
          ((data_in == 2'b01) && soft_reset_1) ||
			 ((data_in == 2'b10) && soft_reset_2))
  state <= DA;
  else
  state <= next_state;
  
  end
  
  always@(state, pkt_valid, data_in, fifo_empty_0, fifo_empty_1, fifo_empty_2, fifo_full, parity_done, low_packet_valid)
  begin
  
  case(state)
  DA : begin
	     if((pkt_valid && (data_in == 2'b00) && fifo_empty_0) || //pkt_valid, data_in, fifo_empty_0, fifo_empty_1, fifo_empty_2
	        (pkt_valid && (data_in == 2'b01) && fifo_empty_1) ||
		    (pkt_valid && (data_in == 2'b10) && fifo_empty_2))
         next_state = LFD;
		 else if((pkt_valid && (data_in == 2'b00) && !fifo_empty_0) ||
	             (pkt_valid && (data_in == 2'b01) && !fifo_empty_1) ||
		         (pkt_valid && (data_in == 2'b10) && !fifo_empty_2))
		 next_state = WTE;
         else
         next_state = DA;
	   end
  
  LFD: next_state = LD;
  
  LD : begin
	     if(!fifo_full && !pkt_valid)
		 next_state = LP;
		 else if(fifo_full)
		 next_state = FFS;
		 else
		 next_state = LD;
       end
	   
  LP : next_state = CPE;
  
  FFS: begin
         if(!fifo_full)
		 next_state = LAF;
		 else
		 next_state = FFS;
	   end
  
  LAF: begin
         if(parity_done)
	     next_state = DA;
	     else if(!parity_done && low_packet_valid)
	     next_state = LP;
	     else if(!parity_done && !low_packet_valid)
	     next_state = LD;
	   end
  
  WTE: begin
         if(((data_in == 2'b00) && fifo_empty_0) ||
	        ((data_in == 2'b01) && fifo_empty_1) ||
		    ((data_in == 2'b10) && fifo_empty_2))
	     next_state = LFD;
		 else
		 next_state = WTE;
	   end
  
  CPE: begin
         if(fifo_full)
	     next_state = FFS;
		 else
		 next_state = DA;
       end
  
  default: next_state = DA;
  endcase  
		
  end

  assign write_enb_reg = ((state == LD) || (state == LP) || (state == LAF)) ? 1'b1 : 1'b0;
  assign detect_add = (state == DA) ? 1'b1 : 1'b0;
  assign ld_state = (state == LD) ? 1'b1 : 1'b0;
  assign laf_state = (state == LAF) ? 1'b1 : 1'b0;
  assign lfd_state = (state == LFD) ? 1'b1 : 1'b0;
  assign full_state = (state == FFS) ? 1'b1 : 1'b0;
  assign rst_int_reg = (state == CPE) ? 1'b1 : 1'b0;
  //assign busy = (state != DA || state != LD) ? 1'b1 : 1'b0;
  //assign busy = state != LD ? 1'b1 : 1'b0;
  assign busy = ((state == LFD) || (state == LP) || (state == FFS) || (state == LAF) || (state == WTE) || (state == CPE)) ? 1'b1 : 1'b0;
  
  endmodule